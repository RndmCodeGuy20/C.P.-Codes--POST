library ieee;
use ieee.std_logic_1164.all;

entity Exp2 is
  port (
    A,B : in std_logic;
    LHS,RHS : out std_logic
  ) ;
end Exp2;